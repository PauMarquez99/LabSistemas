entity Full_Add is

end Full_Add;
