library ieee;
use ieee.std_logic_1164.all;

entity OutputRegister is
  port(O_enb: in std_logic;
    input: in std_logic_vector(3 downto 0);
    Data_O: out std_logic_vector(3 downto 0)
  );
end entity;

architecture log of OutputRegister is

begin
  

end log;
